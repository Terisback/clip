module main

import remimimimi.clip

fn main() {
	println(os.args)
}