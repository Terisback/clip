module clip

fn (app App) parse(args string) ?Matches {
	return none
}
